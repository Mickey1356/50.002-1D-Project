module tile_bitmap (
    input clk,  // clock
    input rst,  // reset
    input enabled,
    input wire [1:0] type,
    input wire [5:0] yline,
    output reg [59:0] bitmap
  );
  
  reg [1:0] rtype;
  reg [5:0] ryline;
  reg [7:0] raddr;

  /* Sequential Logic */
  always @(posedge clk) begin
    if (enabled)
      rtype <= type;
      ryline <= yline;
      raddr <= {type, yline};
  end
  
  always @(raddr) begin
    if (enabled)
      case (raddr)
        8'b00000000: bitmap <= 60'b111111111111111111111111111111111111111111111111111111111111;
        8'b00000001: bitmap <= 60'b111111111111111111111111111111111111111111111111111111111111;
        8'b00000010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00000011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00000100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00000101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00000110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00000111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00001111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00010111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00011111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00100111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00101111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110010: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110011: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110100: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110101: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110110: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00110111: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00111000: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00111001: bitmap <= 60'b110000000000000000000000000000000000000000000000000000000011;
        8'b00111010: bitmap <= 60'b111111111111111111111111111111111111111111111111111111111111;
        8'b00111011: bitmap <= 60'b111111111111111111111111111111111111111111111111111111111111;
        default: bitmap <= 0;
      endcase
  end
  
endmodule
